library verilog;
use verilog.vl_types.all;
entity Fetch_Cycle_tb is
end Fetch_Cycle_tb;
